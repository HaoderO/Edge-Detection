LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY AD7606_DRIVER IS
	PORT
	(
		CLK      	: IN  	STD_LOGIC;                       --时钟75MHz
		BUSY     	: IN  	STD_LOGIC;                       --AD7606开始转换信号
		FIRSTDATA	: IN  	STD_LOGIC;                       --第一个通道输出标志
		INDATA   	: IN  	STD_LOGIC_VECTOR(15 DOWNTO 0);   --16位采样结果
		RESTOUT  	: OUT	STD_LOGIC;                       --AD7606复位信号
		OUTDATA  	: OUT 	STD_LOGIC_VECTOR(15 DOWNTO 0);   --16位采样结果
		ARESS    	: OUT 	STD_LOGIC_VECTOR(3 DOWNTO 0);    --通道
		CONVENT4 	: OUT 	STD_LOGIC;                       --AD7606开始转换信号
		CS       	: OUT 	STD_LOGIC;                       --AD7606下一通道输出信号
		RD       	: OUT 	STD_LOGIC;                       --AD7606下一通道输出信号
		CH_EN    	: OUT 	STD_LOGIC                        --通道数据有效标志
	);
		  
END ENTITY AD7606_DRIVER; 

ARCHITECTURE ART OF AD7606_DRIVER IS
COMPONENT REST IS
PORT
	(
		CLK			: IN 	STD_LOGIC;
		SYS_RET_N	: IN 	STD_LOGIC;
		RSET0		: OUT	STD_LOGIC;
		EN			: OUT	STD_LOGIC
	);
END COMPONENT REST;


COMPONENT CONVENT IS     --控制AD7606开始转换 
PORT
	(
		CLK	    	: IN 	STD_LOGIC;
		EN 	    	: IN    STD_LOGIC;
		FIRSTDATA 	: IN    STD_LOGIC;
		STARTREAD 	: IN	STD_LOGIC;
		ADDRESS   	: IN 	STD_LOGIC_VECTOR(3 DOWNTO 0);
		CONVENT1	: OUT   STD_LOGIC
	);
END COMPONENT CONVENT;
	
	
	
COMPONENT  READ1 IS     --读取AD7606各个通道的采样数据
PORT
	(
		CLK	    	: IN 	STD_LOGIC;
		EN 	    	: IN    STD_LOGIC;
		CONVENT1  	: IN    STD_LOGIC;
		BUSY      	: IN	STD_LOGIC;
		FIRSTDATA 	: IN	STD_LOGIC;
		INDATA	 	: IN 	STD_LOGIC_VECTOR(15 DOWNTO 0);
		RD    	 	: OUT   STD_LOGIC;
		OUTDATA	 	: OUT	STD_LOGIC_VECTOR(15 DOWNTO 0);
		STARTREAD1	: OUT 	STD_LOGIC;
		ADDRESS	 	: OUT   STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT READ1;


COMPONENT  HIGN IS    --AD7606各个通道数据输出有效
PORT
	(
		CLK			: IN 	STD_LOGIC;
		ARESS		: IN 	STD_LOGIC_VECTOR(3 DOWNTO 0);
		CH_EN		: OUT 	STD_LOGIC
	);
END COMPONENT HIGN;




SIGNAL EN,RSET12,CONVENT12:STD_LOGIC;
SIGNAL CLK1,CLK2      	  :STD_LOGIC;
SIGNAL RESTIN             :STD_LOGIC:='1';
SIGNAL STARTREAD4,CSRD    :STD_LOGIC;
SIGNAL ADDRESS            :STD_LOGIC_VECTOR(3 DOWNTO 0);

BEGIN
U1:REST     PORT MAP(CLK,RESTIN,RESTOUT,EN);
U2:CONVENT  PORT MAP(CLK,EN,FIRSTDATA,STARTREAD4,ADDRESS,CONVENT12);
U3:READ1    PORT MAP(CLK,EN,CONVENT12,BUSY,FIRSTDATA,INDATA,CSRD,OUTDATA,STARTREAD4,ADDRESS);
U5:HIGN     PORT MAP(CLK,ADDRESS,CH_EN);

ARESS<=ADDRESS;
CONVENT4<=CONVENT12;
CS<=CSRD;
RD<=CSRD;

END ARCHITECTURE ART;