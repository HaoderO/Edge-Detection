LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
--此模块的作用是判断AD是否正在输出8个通道数据
--高电平阶段表示AD正输出8个通道数据
ENTITY HIGN IS
	PORT(
			CLK	: IN 	STD_LOGIC;
			ARESS	: IN 	STD_LOGIC_VECTOR(3 DOWNTO 0);
			CH_EN	: OUT STD_LOGIC
			);
END ENTITY HIGN;

ARCHITECTURE ART OF HIGN IS

BEGIN

PROCESS(ARESS,CLK)--判断AD是否正在输出8个通道数据
BEGIN
	IF(CLK'EVENT AND CLK='1')THEN
		IF (ARESS>="0001" AND ARESS<="1000") THEN 
			CH_EN<='1';    
		ELSE
			CH_EN<='0'; 
		END IF;			
	END IF;
END PROCESS;
	
END ARCHITECTURE ART;