LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY FPGAWR_DSPRE_CTRL IS
PORT (
        SYS_CLK     : IN     STD_LOGIC;--75MHz
        XA          : IN     STD_LOGIC_VECTOR(11 DOWNTO 0); --12位地址总线
        XZCS_7      : IN     STD_LOGIC := '1';              --ZONE7片选使能
        XRD         : IN     STD_LOGIC := '1';              --DSP读使能
 
        WREN_A      : BUFFER STD_LOGIC := '0';              --RAM_A读使能
        RDEN_A      : BUFFER STD_LOGIC := '0';              --RAM_A写使能
        ADDRESS_A   : BUFFER STD_LOGIC_VECTOR(11 DOWNTO 0) := "000000000000";--FPGA写数据地址
        ADDRESS_CH  : IN     STD_LOGIC_VECTOR(3 DOWNTO 0);  --AD通道序号
        VALID_FLAG  : IN     STD_LOGIC                      --AD数据有效标志
    );
END ENTITY;

ARCHITECTURE A OF FPGAWR_DSPRE_CTRL IS

SIGNAL ADDR_FPGAWR  : STD_LOGIC_VECTOR(11 DOWNTO 0) := "000000000000";--FPGA写地址计数信号
SIGNAL CH_CNT       : STD_LOGIC_VECTOR(11 DOWNTO 0) := "000000000000";--FPGA写地址计数的基数信号

BEGIN

READ_EN : PROCESS(XRD,XZCS_7)           --RAM_A读使能判断
BEGIN
    IF((XZCS_7='0')AND(XRD='0')) THEN
	RDEN_A <= '1';
    ELSE
	RDEN_A <= '0';
    END IF;
END PROCESS;

WRITE_EN : PROCESS(VALID_FLAG,RDEN_A)   --RAM_A写使能判断
BEGIN
	IF((VALID_FLAG='1')AND(RDEN_A='0')) THEN
		WREN_A <= '1';
    ELSE        
        WREN_A <= '0';
	END IF;
END PROCESS;

ADDRESS_SWAP : PROCESS(XRD,XZCS_7)      --RAM_A读写地址切换
BEGIN
    IF((XZCS_7='0')AND(XRD='0')) THEN
        ADDRESS_A <= XA;                --DSP读数据时地址由DSP提供
    ELSE
        ADDRESS_A <= ADDR_FPGAWR;       --FPGA写数据时地址由FPGA提供
    END IF;
END PROCESS;

PROCESS(VALID_FLAG,CH_CNT)                     --生成FPGA写地址地址基数
BEGIN
    IF(VALID_FLAG'EVENT AND VALID_FLAG='1') THEN
        IF(CH_CNT="011111111000") THEN
            CH_CNT <= "000000000000"; 
	    ELSE
            CH_CNT <= CH_CNT  + "000000001000";--VALID_FLAG上升沿地址基数加8
	    END IF;
    END IF;
END PROCESS;

ADDRESS_CNT : PROCESS(WREN_A,ADDR_FPGAWR)--生成FPGA写数据地址(0~2047)
BEGIN
    IF(WREN_A='1') THEN
	    IF(ADDR_FPGAWR="011111111111") THEN
	    	ADDR_FPGAWR <= "000000000000";
	    ELSE
	    	ADDR_FPGAWR <= CH_CNT + (ADDRESS_CH-"0001");--FPGA写地址=地址基数+AD数据通道序号
	    END IF;
    END IF;
END PROCESS;

END A;