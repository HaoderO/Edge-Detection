LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DATABUS_SWAP_tb IS 
END DATABUS_SWAP_tb;

ARCHITECTURE TESTBENCH_ARCH OF DATABUS_SWAP_tb IS

COMPONENT DATABUS_SWAP
PORT (
--        SYS_CLK     : IN     STD_LOGIC;
        XRD         : IN     STD_LOGIC;
        XWE         : IN     STD_LOGIC;
		XD          : INOUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		Q_A         : IN     STD_LOGIC_VECTOR(15 DOWNTO 0);
		DATA_B      : OUT    STD_LOGIC_VECTOR(15 DOWNTO 0)
    );
END COMPONENT;

--COMPONENT DA_DATA
--PORT(
--        SYS_CLK     : IN     STD_LOGIC;
--        Q_DATA      : BUFFER STD_LOGIC_VECTOR(15 DOWNTO 0) := "0000000000000000"
--    );
--END COMPONENT;


SIGNAL SYS_CLK      : STD_LOGIC;
SIGNAL XRD          : STD_LOGIC := '0';
SIGNAL XWE          : STD_LOGIC := '0';
SIGNAL XD           : STD_LOGIC_VECTOR(15 DOWNTO 0) := "0000000000000000";
SIGNAL Q_A          : STD_LOGIC_VECTOR(15 DOWNTO 0) := "0000000000000000";
SIGNAL DATA_B       : STD_LOGIC_VECTOR(15 DOWNTO 0) := "0000000000000000";
SIGNAL Q_DATA       : STD_LOGIC_VECTOR(15 DOWNTO 0) := "0000000000000000";

--SIGNAL XD_CHANGE    : STD_LOGIC := '0';

CONSTANT CLK_PERIOD : TIME := 40 NS;

BEGIN

INSTANT1: DATABUS_SWAP PORT MAP
	(
--        SYS_CLK     =>SYS_CLK   , 
		XRD         =>XRD       ,   
		XWE      	=>XWE       ,    
		XD       	=>XD        ,    
        Q_A      	=>Q_A       ,   
        DATA_B      =>DATA_B   
	);

CLK_IN: PROCESS
BEGIN
    SYS_CLK <= '0';
	WAIT FOR CLK_PERIOD/2;
    SYS_CLK <= '1';
	WAIT FOR CLK_PERIOD/2;
END PROCESS;

PROCESS
BEGIN
    XRD <= '1';
    XWE <= '0';
	WAIT FOR CLK_PERIOD*16;
    XRD <= '0';
    XWE <= '1';
	WAIT FOR CLK_PERIOD*16;
END PROCESS;

PROCESS(SYS_CLK)
BEGIN
    IF((XRD='1')AND(XWE='0')) THEN 
    ELSIF(SYS_CLK'EVENT AND SYS_CLK='0') THEN 
        IF(Q_A="0000000000001111") THEN
            Q_A <= "0000000000000000";
        ELSE
            Q_A <= Q_A + '1';
        END IF;
    END IF;
END PROCESS;

PROCESS(XRD,XWE)
BEGIN
    IF((XRD='0')OR(XWE='1')) THEN 
--    ELSIF(SYS_CLK'EVENT AND SYS_CLK='0') THEN 
    	IF(Q_DATA="0000000000100000") THEN
            Q_DATA <= "0000000000000000";
    	ELSE
           	Q_DATA <= Q_DATA + '1';
    	END IF;
    END IF;
END PROCESS;

PROCESS(XRD,XWE)
BEGIN
    IF((XRD='1')AND(XWE='0')) THEN 
        XD <= Q_DATA;
    ELSE
        XD <= "ZZZZZZZZZZZZZZZZ";
    END IF; 
END PROCESS;

END TESTBENCH_ARCH;