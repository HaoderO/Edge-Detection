LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_SIGNED.ALL;
ENTITY REST IS
	PORT(
			CLK			: IN 	STD_LOGIC;
			SYS_RET_N	: IN 	STD_LOGIC;
			RSET0		: OUT 	STD_LOGIC;
			EN			: OUT 	STD_LOGIC
		);
END ENTITY REST;

ARCHITECTURE ART OF REST IS

SIGNAL CQI:	STD_LOGIC_VECTOR(4 DOWNTO 0) :="00000";   --定义保存计数值的信号CQI

BEGIN

PROCESS(SYS_RET_N,CLK)			--计数信号计数
BEGIN
	IF (SYS_RET_N ='0') THEN 
		CQI<=	"00000";    
	ELSIF( CLK'EVENT AND CLK='1')THEN 
		IF (CQI ="11111") THEN 
			CQI <=CQI;
		ELSE
			CQI<=	CQI + '1';
		END IF;			
	END IF;
END PROCESS;
	
PROCESS(SYS_RET_N,CLK,CQI) 		--输出给AD7606复位信号
BEGIN
	IF SYS_RET_N ='0' THEN 
		RSET0<='0';    
	ELSIF( CLK'EVENT AND CLK='1')THEN 
		IF (CQI ="10000") THEN 
			RSET0<='1';  
		ELSIF(CQI="11011")THEN
			RSET0<='0';
		END IF;
	END IF;
END PROCESS;
	
	
PROCESS(SYS_RET_N,CLK,CQI) 		--使能信号输出
BEGIN
	IF SYS_RET_N ='0' THEN 
		EN<='0';    
	ELSIF( CLK'EVENT AND CLK='1')THEN 
		IF CQI ="11110" THEN 
			EN<='1';    
		END IF;
	END IF;
END PROCESS;
	
END ARCHITECTURE ART;