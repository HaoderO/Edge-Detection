LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DSPWR_FPGARE_CTRL IS
PORT (
        SYS_CLK     : IN     STD_LOGIC;						--75MHz
        XA          : IN     STD_LOGIC_VECTOR(11 DOWNTO 0);	--12位地址总线
        XZCS_7      : IN     STD_LOGIC := '1';				--ZONE7片选使能
        XWE         : IN     STD_LOGIC := '1';				--DSP写使能

        RDEN_B      : BUFFER STD_LOGIC := '1';				--RAM_B读使能
        WREN_B      : BUFFER STD_LOGIC := '0';				--RAM_B写使能
		ADDRESS_B   : BUFFER STD_LOGIC_VECTOR(11 DOWNTO 0)	--FPGA读数据地址
    );
END ENTITY;

ARCHITECTURE A OF DSPWR_FPGARE_CTRL IS

SIGNAL ADDR_FPGARE  : STD_LOGIC_VECTOR(11 DOWNTO 0) := "100000000000"; --FPGA读地址计数信号

BEGIN

WRITE_EN : PROCESS(XWE,XZCS_7)		--RAM_B写使能判断
BEGIN
	IF((XZCS_7='0')AND(XWE='0')) THEN
		WREN_B <= '1';
	ELSE
		WREN_B <= '0';
	END IF;
END PROCESS;

READ_EN : PROCESS(WREN_B,XWE)		--RAM_B读使能判断
BEGIN
	IF((WREN_B='0')AND(XWE='1')) THEN
		RDEN_B <= '1';
	ELSE
		RDEN_B <= '0';
	END IF;
END PROCESS;

ADDRESS_SWAP : PROCESS(XWE,XZCS_7)	--RAM_B读写地址切换
BEGIN
	IF((XZCS_7='0')AND(XWE='0')) THEN
		ADDRESS_B <= XA;			--DSP写数据时地址由DSP提供
	ELSE
		ADDRESS_B <= ADDR_FPGARE;	--FPGA读数据时地址由FPGA提供
	END IF;
END PROCESS;

ADDRESS_CNT : PROCESS(WREN_B)		--生成FPGA读数据地址(2048~4095)
BEGIN
    IF(WREN_B'EVENT AND WREN_B='0') THEN
		IF(ADDR_FPGARE="111111111111") THEN
			ADDR_FPGARE <= "100000000000";
		ELSE
			ADDR_FPGARE <= ADDR_FPGARE + '1';
		END IF;
	END IF;
END PROCESS;

END A;