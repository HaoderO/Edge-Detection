LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_SIGNED.ALL;

ENTITY CONVENT IS
	PORT(
			CLK	    : IN 	STD_LOGIC;
			EN 	    : IN    STD_LOGIC;
			FIRSTDATA : IN    STD_LOGIC;
			STARTREAD : IN		STD_LOGIC;
			ADDRESS   : IN 	STD_LOGIC_VECTOR(3 DOWNTO 0);
			CONVENT1	 : OUT   STD_LOGIC);
			
END ENTITY CONVENT;

--该模块读取通道数，输出CONVENT信号，开始AD7606转换
ARCHITECTURE ART OF CONVENT IS

SIGNAL CQI:	STD_LOGIC_VECTOR(3 DOWNTO 0) :="0000"; 

BEGIN
	
PROCESS(EN,CLK) --上电后计数，当计数到1001，CONVENT输出高电平，AD7606开始转换
BEGIN 
	IF(CLK'EVENT AND CLK='1')THEN 
		IF (EN='0')THEN
			CQI<="0000";
		ELSIF (CQI="1001")THEN
			CQI<=CQI;
		ELSE 
			CQI<=	CQI + '1';
		END IF;
	END IF;
END PROCESS;
	
PROCESS(EN,CLK) --根据时钟CLK、通道数ADDRESS控制CONVENT
BEGIN 
	IF( CLK'EVENT AND CLK='1')THEN 
		IF (EN='1') THEN 
			IF(CQI="0011")THEN
				CONVENT1<='1';
			ELSIF(ADDRESS="1000"AND STARTREAD='1')THEN
				CONVENT1<='1';
			ELSIF(ADDRESS="0100")THEN
				CONVENT1<='0';
			END IF;
		ELSE 
			CONVENT1<='0';
		END IF;
	END IF;
END PROCESS;	

END ARCHITECTURE ART;